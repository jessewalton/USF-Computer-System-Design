// Module Name:    ac97commands 

`timescale 1ns / 1ps

module ac97commands (clock, ready, command_address, command_data,
   command_valid, volume, source);

   input clock;
   input ready;
   output [7:0] command_address;
   output [15:0] command_data;
   output command_valid;
   input [4:0] volume;
   input [2:0] source;

   reg [23:0] command;
   reg command_valid;

   reg [3:0] state;

   assign command_address = command[23:16];
   assign command_data = command[15:0];

   wire [4:0] vol;
   assign vol = 31-volume;  // convert to attenuation
   
   initial begin
      command <= 4'h0;
      // synthesis attribute init of command is "0";
      command_valid <= 1'b0;
      // synthesis attribute init of command_valid is "0";
      //done <= 1'b0;

      // synthesis attribute init of old_ready is "0";
      state <= 16'h0000;
      // synthesis attribute init of state is "0000";
   end

   always @(posedge clock) begin
      if (ready) state <= state+1;

      case (state)
         4'h0: // Read ID
         begin
            command <= 24'h80_0000;
            command_valid <= 1'b1;
         end
         4'h1: // Read ID
            command <= 24'h80_0000;
         4'h3: // headphone volume
            command <= { 8'h04, 3'b000, vol, 3'b000, vol };
         4'h5: // PCM volume
            command <= 24'h18_0808;
         4'h6: // Record source select
            command <= { 8'h1A, 5'b00000, source, 5'b00000, source};
         4'h7: // Record gain = max
            command <= 24'h1C_0F0F;
         4'h9: // set +20db mic gain
            command <= 24'h0E_8048;
         4'hA: // Set beep volume
            command <= 24'h0A_0000;
         4'hB: // PCM out bypass mix1
            command <= 24'h20_8000;
         default:
            command <= 24'h80_0000;
      endcase // case(state)
   
   end // always @ (posedge clock)
endmodule // ac97commands
